package pkg;

import uvm_pkg::*;
`include "uvm_macros.svh"

`include "seq_item.sv"
`include "reg_pkg.sv"
`include "reg2axi_adapter.sv"
`include "sequencer.sv"


`include "driver.sv"
`include "moniter.sv"
`include "agent.sv"
`include "env.sv"
`include "base_seq.sv"
//`include "base_test.sv"
endpackage
